interface siso_if(input logic clk);
  logic rst;
  bit din;
  bit dout;

endinterface
