package my_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "packet.sv"
`include "sequencer.sv"
`include "sequence.sv"

`include "driver.sv"
`include "monitor.sv"
`include "scoreboard.sv"
`include "coverage.sv"
`include "agent.sv"
`include "env.sv"
`include "test.sv"

endpackage : my_pkg



